LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;
--****2015210078 �ſ�****
--LED����ˢ��
--�ڲ����Ԥ��ͼƬ���ⲿ����
--����ʱ�ӽ����л�
--����PWMģ���������
--********2017.11********
ENTITY LEDRefresh IS
    GENERIC (IMGNUM : INTEGER := 6);
	PORT(Rollclock:IN STD_LOGIC;                        --ѭ��ʱ��(����ͼƬƽ��)
        PWMclock:IN STD_LOGIC;                          --PWM����Ƶ��(ӦΪ���������Ƶ�ʵ�256�����ƻ�256KHz����)
        Switchclock:IN STD_LOGIC;                       --��ɨ��Ƶ��(Ӧ����ˢ���ʵ�8�����ƻ�160Hz����)
		LEDEnable:IN STD_LOGIC;                         --����ʹ��
        reset:IN STD_LOGIC;                             --��λ
		luma:IN INTEGER  RANGE 0 TO 255;                --����(ֱ�������PWM��Ϊռ�ձ�)
		DataSel: IN INTEGER  RANGE 0 TO IMGNUM-1;       --ͼ��ѡ��
		Lineout: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);      --����п��ź�
        Columnout: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));  --����п��ź�
END LEDRefresh;
ARCHITECTURE LEDRefresher OF LEDRefresh IS
	COMPONENT PWM
        GENERIC (n : INTEGER := 255);
        PORT(PWMclock:IN STD_LOGIC;     --PWM����Ƶ��(ӦΪ���������Ƶ�ʵ�256��)
		reset:IN STD_LOGIC;             --����
		div:IN INTEGER  RANGE 0 TO n;   --ռ�ձ�0-255
		output:OUT STD_LOGIC);          --���
	END COMPONENT;
    COMPONENT RollGate IS
        PORT(Rollclock:IN STD_LOGIC;
            reset:IN STD_LOGIC;
            Enable:IN STD_LOGIC;
            Direction:IN STD_LOGIC;                     --0��1��
            input:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            output:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
    END COMPONENT;
	SIGNAL PwmWave:STD_LOGIC;                               --PWM����ź���
    SIGNAL lcount:INTEGER RANGE 0 TO 7;                     --�м�����
    SIGNAL RollEnable:STD_LOGIC;                            --ѭ��ʹ��
    SIGNAL Direction:STD_LOGIC;                             --ѭ��ʹ��
    SIGNAL ColumnSignal: STD_LOGIC_VECTOR(15 DOWNTO 0);     --����п��ź�
                        --ͼƬ��6             ����8      ����16
    TYPE IMGS IS ARRAY (IMGNUM-1 DOWNTO 0,7 DOWNTO 0,15 DOWNTO 0) OF STD_LOGIC;
    --IMG����Գ�
    CONSTANT Data:IMGS:=
                (	--5
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('0','0','0','0','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','0','0','0','0','0' , '0','0','1','0','0','1','0','0'),
                        ('0','0','1','0','0','1','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','1','0','0','1','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','1','1','1','1','1','1','0' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '1','1','1','1','1','1','1','1'),
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0')
                    ),
                    --4
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '1','1','1','1','1','1','1','1'),
                        ('1','1','1','1','1','1','1','1' , '1','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1')
                    ),
                    --3
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('0','0','0','0','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','1','0','0','0','0','1','0' , '0','0','0','1','1','0','0','0'),
                        ('1','0','0','0','0','0','0','1' , '0','0','0','1','1','0','0','0'),
                        ('0','1','1','1','1','1','1','0' , '0','0','0','0','0','0','0','0'),
                        ('1','1','0','0','0','1','1','0' , '0','0','0','0','0','0','0','0'),
                        ('0','1','0','0','0','0','1','0' , '0','1','0','0','0','0','1','0'),
                        ('1','0','1','0','0','1','0','1' , '1','0','1','0','0','1','0','1'),
                        ('0','1','0','0','0','0','1','0' , '0','1','0','0','0','0','1','0' )
                    ),
                    --2ͣ��
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('0','0','0','0','0','0','0','0' , '1','0','0','0','0','0','0','1'),
                        ('0','0','0','0','0','0','0','0' , '0','1','0','0','0','0','1','0'),
                        ('0','0','0','0','0','0','0','0' , '0','0','1','0','0','1','0','0'),
                        ('0','0','0','0','0','0','0','0' , '0','0','0','1','1','0','0','0'),
                        ('0','0','0','0','0','0','0','0' , '0','0','0','1','1','0','0','0'),
                        ('0','0','0','0','0','0','0','0' , '0','0','1','0','0','1','0','0'),
                        ('0','0','0','0','0','0','0','0' , '0','1','0','0','0','0','1','0'),
                        ('0','0','0','0','0','0','0','0' , '1','0','0','0','0','0','0','1')
                    ),
                    --1��ͷ
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('0','0','0','0','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','0','1','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','0','0','1','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','0','0','0','1','0' , '0','0','0','0','0','0','0','0'),
                        ('0','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','0','0','0','1','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','0','0','1','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','0','1','0','0','0' , '0','0','0','0','0','0','0','0')
                    ),
                    --0��ͷ
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('0','0','0','0','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','1','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','1','0','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','1','0','0','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','0' , '0','0','0','0','0','0','0','0'),
                        ('0','1','0','0','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','1','0','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','1','0','0','0','0' , '0','0','0','0','0','0','0','0')
                    )
                );
BEGIN
	PWMGen: PWM PORT MAP (PWMclock=>PWMclock,reset=>reset,div=>luma,output=>PwmWave);
    RedLEDP : RollGate PORT MAP (Rollclock=>Rollclock,reset=>reset,Enable=>RollEnable,
    Direction=>Direction,input=>ColumnSignal(7 DOWNTO 0),output=>Columnout(7 DOWNTO 0));
    GreenLEDP : RollGate PORT MAP (Rollclock=>Rollclock,reset=>reset,Enable=>RollEnable,
    Direction=>Direction,input=>ColumnSignal(15 DOWNTO 8),output=>Columnout(15 DOWNTO 8));
	PROCESS(Rollclock,Switchclock,lcount,DataSel,PwmWave,LEDEnable,reset)
	BEGIN
		IF(LEDEnable='0' OR reset='1')THEN
			ColumnSignal<=std_logic_vector(to_unsigned(0, 16));
            Lineout<="11111111";
            RollEnable <= '0';
            Direction <= '1';
		ELSE
            --LED��ˢ�¼���
            IF(Switchclock'event AND Switchclock='0')THEN
                lcount<=lcount+1;
            END IF;
            --LED��ѡ ѡ�е�һ�����źŵ͵�λ,δѡ�е������źŸߵ�λ
            Lineout <= NOT TO_STDLOGICVECTOR("00000001" SLL lcount);
            --��ʾһ��
            IF(DataSel = 0)THEN     --��תͼƬ
                RollEnable <= '1';  --ͼƬ����ʹ��
                Direction <= '0';   --���ù�������
            ELSIF(DataSel = 1)THEN  --��תͼƬ
                RollEnable <= '1';
                Direction <= '1';
            ELSE                    --����ͼƬ
                RollEnable <= '0';  --����ͼƬ����
                Direction <= '1';   --���ù�������(�˴���������)
            END IF;
            FOR c IN 0 TO 15 LOOP
                IF Data(DataSel,lcount,c)='1' THEN                   
                    ColumnSignal(c) <= PwmWave;--ѡ�е�һ�����ź�PWM��λ
                ELSE
                    ColumnSignal(c) <= '0';    --δѡ�е�һ�����źŵ͵�λ
                END IF;                                     
            END LOOP;                                     
		END IF;
	END PROCESS;
END LEDRefresher;