LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;
--------------------------------
--LED����ˢ��
--�ڲ����Ԥ��ͼƬ���ⲿ����
--����ʱ�ӽ����л�
--����PWMģ���������
--
--------------------------------

ENTITY LEDRefresh IS
    GENERIC (IMGNUM : INTEGER := 6);
	PORT(Rollclock:IN STD_LOGIC;                        --ѭ��ʱ��
        PWMclock:IN STD_LOGIC;                          --PWM����Ƶ��(ӦΪ���������Ƶ�ʵ�256�����ƻ�256KHz����)
        Switchclock:IN STD_LOGIC;                       --��ɨ��Ƶ��(Ӧ����ˢ���ʵ�8�����ƻ�160Hz����)
		LEDEnable:IN STD_LOGIC;                         --����ʹ��
        reset:IN STD_LOGIC;                             --��λ
		luma:IN INTEGER  RANGE 0 TO 255;                --����(ֱ�������PWM��Ϊռ�ձ�)
		DataSel: IN INTEGER  RANGE 0 TO IMGNUM-1;       --ͼ��ѡ��
		Lineout: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);      --����п��ź�
        Columnout: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));  --����п��ź�
END LEDRefresh;
ARCHITECTURE LEDRefresher OF LEDRefresh IS
	COMPONENT PWM
		PORT(PWMclock:IN STD_LOGIC;
		reset:IN STD_LOGIC;
		div:IN INTEGER  RANGE 0 TO 255;
		output:OUT STD_LOGIC);
	END COMPONENT;
	SIGNAL PwmWave:STD_LOGIC;               --PWM����ź���
    SIGNAL lcount:INTEGER RANGE 0 TO 7;     --�м�����
                        --ͼƬ��    ����        ����
    --TYPE LINEP IS ARRAY (15 DOWNTO 0) OF STD_LOGIC;
    --TYPE IMG IS ARRAY (7 DOWNTO 0) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
    TYPE IMGS IS ARRAY (IMGNUM-1 DOWNTO 0,7 DOWNTO 0) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
    --TYPE IMGS IS ARRAY (IMGNUM-1 DOWNTO 0,7 DOWNTO 0,15 DOWNTO 0) OF STD_LOGIC;
    --IMG����Գ�
    SIGNAL Data:IMGS;
BEGIN
	PWMGen: PWM PORT MAP (PWMclock=>PWMclock,reset=>reset,div=>luma,output=>PwmWave);
	PROCESS(Rollclock,Switchclock,lcount,DataSel,PwmWave,LEDEnable,reset,Data)
	BEGIN
		IF(LEDEnable='0' OR reset='1')THEN
			Columnout<=std_logic_vector(to_unsigned(0, 16));
            Lineout<="11111111";
            Data<=
                (	--5
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '1','0','1','0','1','0','1','0'),
                        ('0','1','0','1','0','1','0','1' , '1','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1')
                    ),
                    --4
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('0','1','0','1','0','1','0','1' , '1','0','1','0','1','0','1','0'),
                        ('0','1','0','1','0','1','0','1' , '1','0','1','0','1','0','1','0'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1')
                    ),
                    --3
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','1' , '0','0','0','0','0','0','0','0'),
                        ('0','1','0','1','0','1','0','1' , '1','1','1','1','1','1','1','1'),
                        ('1','1','1','1','1','1','1','1' , '1','0','1','0','1','0','1','0'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','0','0' , '1','1','1','1','1','1','1','1')
                    ),
                    --2ͣ��
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('0','0','0','0','0','0','0','0' , '1','0','0','0','0','0','0','1'),
                        ('0','0','0','0','0','0','0','0' , '0','1','0','0','0','0','1','0'),
                        ('0','0','0','0','0','0','0','0' , '0','0','1','0','0','1','0','0'),
                        ('0','0','0','0','0','0','0','0' , '0','0','0','1','1','0','0','0'),
                        ('0','0','0','0','0','0','0','0' , '0','0','0','1','1','0','0','0'),
                        ('0','0','0','0','0','0','0','0' , '0','0','1','0','0','1','0','0'),
                        ('0','0','0','0','0','0','0','0' , '0','1','0','0','0','0','1','0'),
                        ('0','0','0','0','0','0','0','0' , '1','0','0','0','0','0','0','1')
                    ),
                    --1��ͷ
                    (--  15   14  13  12  11  10  9   8     7   6   5   4   3   2   1   0
                        ('0','0','0','0','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','0','1','0','0','0' , '0','0','0','0','1','0','0','0'),
                        ('0','0','0','0','0','1','0','0' , '0','0','0','0','0','1','0','0'),
                        ('0','0','0','0','0','0','1','0' , '0','0','0','0','0','0','1','0'),
                        ('0','1','1','1','1','1','1','1' , '0','1','1','1','1','1','1','1'),
                        ('0','0','0','0','0','0','1','0' , '0','0','0','0','0','0','1','0'),
                        ('0','0','0','0','0','1','0','0' , '0','0','0','0','0','1','0','0'),
                        ('0','0','0','0','1','0','0','0' , '0','0','0','0','1','0','0','0')
                    ),
                    --0��ͷ
                    (
                        ('0','0','0','0','0','0','0','0' , '0','0','0','0','0','0','0','0'),
                        ('0','0','0','1','0','0','0','0' , '0','0','0','1','0','0','0','0'),
                        ('0','0','1','0','0','0','0','0' , '0','0','1','0','0','0','0','0'),
                        ('0','1','0','0','0','0','0','0' , '0','1','0','0','0','0','0','0'),
                        ('1','1','1','1','1','1','1','0' , '1','1','1','1','1','1','1','0'),
                        ('0','1','0','0','0','0','0','0' , '0','1','0','0','0','0','0','0'),
                        ('0','0','1','0','0','0','0','0' , '0','0','1','0','0','0','0','0'),
                        ('0','0','0','1','0','0','0','0' , '0','0','0','1','0','0','0','0')
                    )
                );
		ELSE
            --����
            IF(Switchclock'event AND Switchclock='0')THEN
                --ѡ��һ��
                lcount<=lcount+1;
            END IF;
            Lineout <= NOT TO_STDLOGICVECTOR("00000001" SLL lcount);--ѡ�е�һ�����źŵ͵�λ,δѡ�е������źŸߵ�λ
            --��ʾһ��
            
            --ѭ��
            IF(Rollclock'event AND Rollclock='0')THEN
                FOR l IN 0 TO 7 LOOP
                    Data(0,l) <= TO_STDLOGICVECTOR(TO_BITVECTOR(Data(DataSel,l)) ROL 1);
                    Data(1,l) <= TO_STDLOGICVECTOR(TO_BITVECTOR(Data(DataSel,l)) ROR 1);
                END LOOP; 
            END IF;
            
            FOR c IN 0 TO 15 LOOP
                IF Data(DataSel,lcount)(c)='1' THEN                   
                    Columnout(c) <= PwmWave;--ѡ�е�һ�����ź�PWM��λ
                ELSE
                    Columnout(c) <= '0';    --δѡ�е�һ�����źŵ͵�λ
                END IF;                                     
            END LOOP;                                     
		END IF;
	END PROCESS;
END LEDRefresher;